module KAN(
    input wire clk,
    input wire rst,
    input wire [31:0] x1,
    input wire [31:0] x2,
    output wire [31:0] y
);

// Intermediate signals
wire [31:0] layer0_out_0;
wire [31:0] layer0_out_1;
wire [31:0] layer0_out_2;
wire [31:0] layer1_out_0;
wire [31:0] layer1_out_1;
wire [31:0] layer1_out_2;
wire [31:0] layer2_out;

reg [7:0] layers_0_base_weight_0;
reg [7:0] layers_0_base_weight_1;
reg [7:0] layers_0_base_weight_2;
reg [7:0] layers_0_base_weight_3;
reg [7:0] layers_0_base_weight_4;
reg [7:0] layers_0_base_weight_5;
reg [7:0] layers_0_spline_scaler_0;
reg [7:0] layers_0_spline_scaler_1;
reg [7:0] layers_0_spline_scaler_2;
reg [7:0] layers_0_spline_scaler_3;
reg [7:0] layers_0_spline_scaler_4;
reg [7:0] layers_0_spline_scaler_5;
reg [7:0] layers_0_spline_weight_0;
reg [7:0] layers_0_spline_weight_1;
reg [7:0] layers_0_spline_weight_2;
reg [7:0] layers_0_spline_weight_3;
reg [7:0] layers_0_spline_weight_4;
reg [7:0] layers_0_spline_weight_5;
reg [7:0] layers_0_spline_weight_6;
reg [7:0] layers_0_spline_weight_7;
reg [7:0] layers_0_spline_weight_8;
reg [7:0] layers_0_spline_weight_9;
reg [7:0] layers_0_spline_weight_10;
reg [7:0] layers_0_spline_weight_11;
reg [7:0] layers_0_spline_weight_12;
reg [7:0] layers_0_spline_weight_13;
reg [7:0] layers_0_spline_weight_14;
reg [7:0] layers_0_spline_weight_15;
reg [7:0] layers_0_spline_weight_16;
reg [7:0] layers_0_spline_weight_17;
reg [7:0] layers_0_spline_weight_18;
reg [7:0] layers_0_spline_weight_19;
reg [7:0] layers_0_spline_weight_20;
reg [7:0] layers_0_spline_weight_21;
reg [7:0] layers_0_spline_weight_22;
reg [7:0] layers_0_spline_weight_23;
reg [7:0] layers_0_spline_weight_24;
reg [7:0] layers_0_spline_weight_25;
reg [7:0] layers_0_spline_weight_26;
reg [7:0] layers_0_spline_weight_27;
reg [7:0] layers_0_spline_weight_28;
reg [7:0] layers_0_spline_weight_29;
reg [7:0] layers_0_spline_weight_30;
reg [7:0] layers_0_spline_weight_31;
reg [7:0] layers_0_spline_weight_32;
reg [7:0] layers_0_spline_weight_33;
reg [7:0] layers_0_spline_weight_34;
reg [7:0] layers_0_spline_weight_35;
reg [7:0] layers_0_spline_weight_36;
reg [7:0] layers_0_spline_weight_37;
reg [7:0] layers_0_spline_weight_38;
reg [7:0] layers_0_spline_weight_39;
reg [7:0] layers_0_spline_weight_40;
reg [7:0] layers_0_spline_weight_41;
reg [7:0] layers_0_spline_weight_42;
reg [7:0] layers_0_spline_weight_43;
reg [7:0] layers_0_spline_weight_44;
reg [7:0] layers_0_spline_weight_45;
reg [7:0] layers_0_spline_weight_46;
reg [7:0] layers_0_spline_weight_47;
reg [7:0] layers_1_base_weight_0;
reg [7:0] layers_1_base_weight_1;
reg [7:0] layers_1_base_weight_2;
reg [7:0] layers_1_base_weight_3;
reg [7:0] layers_1_base_weight_4;
reg [7:0] layers_1_base_weight_5;
reg [7:0] layers_1_base_weight_6;
reg [7:0] layers_1_base_weight_7;
reg [7:0] layers_1_base_weight_8;
reg [7:0] layers_1_spline_scaler_0;
reg [7:0] layers_1_spline_scaler_1;
reg [7:0] layers_1_spline_scaler_2;
reg [7:0] layers_1_spline_scaler_3;
reg [7:0] layers_1_spline_scaler_4;
reg [7:0] layers_1_spline_scaler_5;
reg [7:0] layers_1_spline_scaler_6;
reg [7:0] layers_1_spline_scaler_7;
reg [7:0] layers_1_spline_scaler_8;
reg [7:0] layers_1_spline_weight_0;
reg [7:0] layers_1_spline_weight_1;
reg [7:0] layers_1_spline_weight_2;
reg [7:0] layers_1_spline_weight_3;
reg [7:0] layers_1_spline_weight_4;
reg [7:0] layers_1_spline_weight_5;
reg [7:0] layers_1_spline_weight_6;
reg [7:0] layers_1_spline_weight_7;
reg [7:0] layers_1_spline_weight_8;
reg [7:0] layers_1_spline_weight_9;
reg [7:0] layers_1_spline_weight_10;
reg [7:0] layers_1_spline_weight_11;
reg [7:0] layers_1_spline_weight_12;
reg [7:0] layers_1_spline_weight_13;
reg [7:0] layers_1_spline_weight_14;
reg [7:0] layers_1_spline_weight_15;
reg [7:0] layers_1_spline_weight_16;
reg [7:0] layers_1_spline_weight_17;
reg [7:0] layers_1_spline_weight_18;
reg [7:0] layers_1_spline_weight_19;
reg [7:0] layers_1_spline_weight_20;
reg [7:0] layers_1_spline_weight_21;
reg [7:0] layers_1_spline_weight_22;
reg [7:0] layers_1_spline_weight_23;
reg [7:0] layers_1_spline_weight_24;
reg [7:0] layers_1_spline_weight_25;
reg [7:0] layers_1_spline_weight_26;
reg [7:0] layers_1_spline_weight_27;
reg [7:0] layers_1_spline_weight_28;
reg [7:0] layers_1_spline_weight_29;
reg [7:0] layers_1_spline_weight_30;
reg [7:0] layers_1_spline_weight_31;
reg [7:0] layers_1_spline_weight_32;
reg [7:0] layers_1_spline_weight_33;
reg [7:0] layers_1_spline_weight_34;
reg [7:0] layers_1_spline_weight_35;
reg [7:0] layers_1_spline_weight_36;
reg [7:0] layers_1_spline_weight_37;
reg [7:0] layers_1_spline_weight_38;
reg [7:0] layers_1_spline_weight_39;
reg [7:0] layers_1_spline_weight_40;
reg [7:0] layers_1_spline_weight_41;
reg [7:0] layers_1_spline_weight_42;
reg [7:0] layers_1_spline_weight_43;
reg [7:0] layers_1_spline_weight_44;
reg [7:0] layers_1_spline_weight_45;
reg [7:0] layers_1_spline_weight_46;
reg [7:0] layers_1_spline_weight_47;
reg [7:0] layers_1_spline_weight_48;
reg [7:0] layers_1_spline_weight_49;
reg [7:0] layers_1_spline_weight_50;
reg [7:0] layers_1_spline_weight_51;
reg [7:0] layers_1_spline_weight_52;
reg [7:0] layers_1_spline_weight_53;
reg [7:0] layers_1_spline_weight_54;
reg [7:0] layers_1_spline_weight_55;
reg [7:0] layers_1_spline_weight_56;
reg [7:0] layers_1_spline_weight_57;
reg [7:0] layers_1_spline_weight_58;
reg [7:0] layers_1_spline_weight_59;
reg [7:0] layers_1_spline_weight_60;
reg [7:0] layers_1_spline_weight_61;
reg [7:0] layers_1_spline_weight_62;
reg [7:0] layers_1_spline_weight_63;
reg [7:0] layers_1_spline_weight_64;
reg [7:0] layers_1_spline_weight_65;
reg [7:0] layers_1_spline_weight_66;
reg [7:0] layers_1_spline_weight_67;
reg [7:0] layers_1_spline_weight_68;
reg [7:0] layers_1_spline_weight_69;
reg [7:0] layers_1_spline_weight_70;
reg [7:0] layers_1_spline_weight_71;
reg [7:0] layers_2_base_weight_0;
reg [7:0] layers_2_base_weight_1;
reg [7:0] layers_2_base_weight_2;
reg [7:0] layers_2_spline_scaler_0;
reg [7:0] layers_2_spline_scaler_1;
reg [7:0] layers_2_spline_scaler_2;
reg [7:0] layers_2_spline_weight_0;
reg [7:0] layers_2_spline_weight_1;
reg [7:0] layers_2_spline_weight_2;
reg [7:0] layers_2_spline_weight_3;
reg [7:0] layers_2_spline_weight_4;
reg [7:0] layers_2_spline_weight_5;
reg [7:0] layers_2_spline_weight_6;
reg [7:0] layers_2_spline_weight_7;
reg [7:0] layers_2_spline_weight_8;
reg [7:0] layers_2_spline_weight_9;
reg [7:0] layers_2_spline_weight_10;
reg [7:0] layers_2_spline_weight_11;
reg [7:0] layers_2_spline_weight_12;
reg [7:0] layers_2_spline_weight_13;
reg [7:0] layers_2_spline_weight_14;
reg [7:0] layers_2_spline_weight_15;
reg [7:0] layers_2_spline_weight_16;
reg [7:0] layers_2_spline_weight_17;
reg [7:0] layers_2_spline_weight_18;
reg [7:0] layers_2_spline_weight_19;
reg [7:0] layers_2_spline_weight_20;
reg [7:0] layers_2_spline_weight_21;
reg [7:0] layers_2_spline_weight_22;
reg [7:0] layers_2_spline_weight_23;

initial begin
    layers_0_base_weight_0 = 8'b11111111;
    layers_0_base_weight_1 = 8'b01110010;
    layers_0_base_weight_2 = 8'b11111001;
    layers_0_base_weight_3 = 8'b00000000;
    layers_0_base_weight_4 = 8'b11111110;
    layers_0_base_weight_5 = 8'b11011100;
    layers_0_spline_scaler_0 = 8'b00000000;
    layers_0_spline_scaler_1 = 8'b10010000;
    layers_0_spline_scaler_2 = 8'b10111000;
    layers_0_spline_scaler_3 = 8'b11100101;
    layers_0_spline_scaler_4 = 8'b01110111;
    layers_0_spline_scaler_5 = 8'b11111111;
    layers_0_spline_weight_0 = 8'b10111001;
    layers_0_spline_weight_1 = 8'b11000000;
    layers_0_spline_weight_2 = 8'b11000100;
    layers_0_spline_weight_3 = 8'b10011110;
    layers_0_spline_weight_4 = 8'b11101011;
    layers_0_spline_weight_5 = 8'b11111110;
    layers_0_spline_weight_6 = 8'b01101010;
    layers_0_spline_weight_7 = 8'b10101110;
    layers_0_spline_weight_8 = 8'b10111000;
    layers_0_spline_weight_9 = 8'b10111001;
    layers_0_spline_weight_10 = 8'b10111010;
    layers_0_spline_weight_11 = 8'b10111010;
    layers_0_spline_weight_12 = 8'b10110100;
    layers_0_spline_weight_13 = 8'b10111010;
    layers_0_spline_weight_14 = 8'b10110111;
    layers_0_spline_weight_15 = 8'b10110111;
    layers_0_spline_weight_16 = 8'b10111000;
    layers_0_spline_weight_17 = 8'b10111010;
    layers_0_spline_weight_18 = 8'b10111100;
    layers_0_spline_weight_19 = 8'b10110100;
    layers_0_spline_weight_20 = 8'b10110010;
    layers_0_spline_weight_21 = 8'b10101010;
    layers_0_spline_weight_22 = 8'b10100101;
    layers_0_spline_weight_23 = 8'b10110110;
    layers_0_spline_weight_24 = 8'b10111000;
    layers_0_spline_weight_25 = 8'b10111001;
    layers_0_spline_weight_26 = 8'b10110101;
    layers_0_spline_weight_27 = 8'b10101111;
    layers_0_spline_weight_28 = 8'b10010111;
    layers_0_spline_weight_29 = 8'b10011001;
    layers_0_spline_weight_30 = 8'b10100001;
    layers_0_spline_weight_31 = 8'b10110011;
    layers_0_spline_weight_32 = 8'b10111000;
    layers_0_spline_weight_33 = 8'b10110110;
    layers_0_spline_weight_34 = 8'b10111001;
    layers_0_spline_weight_35 = 8'b11010101;
    layers_0_spline_weight_36 = 8'b11101010;
    layers_0_spline_weight_37 = 8'b11111110;
    layers_0_spline_weight_38 = 8'b11110000;
    layers_0_spline_weight_39 = 8'b10111101;
    layers_0_spline_weight_40 = 8'b10111000;
    layers_0_spline_weight_41 = 8'b10111011;
    layers_0_spline_weight_42 = 8'b10101010;
    layers_0_spline_weight_43 = 8'b10000001;
    layers_0_spline_weight_44 = 8'b00101110;
    layers_0_spline_weight_45 = 8'b00000000;
    layers_0_spline_weight_46 = 8'b01000110;
    layers_0_spline_weight_47 = 8'b10101010;
    layers_1_base_weight_0 = 8'b10101111;
    layers_1_base_weight_1 = 8'b11100110;
    layers_1_base_weight_2 = 8'b10111110;
    layers_1_base_weight_3 = 8'b00101001;
    layers_1_base_weight_4 = 8'b00010000;
    layers_1_base_weight_5 = 8'b01101101;
    layers_1_base_weight_6 = 8'b11111111;
    layers_1_base_weight_7 = 8'b00000010;
    layers_1_base_weight_8 = 8'b00000000;
    layers_1_spline_scaler_0 = 8'b10011001;
    layers_1_spline_scaler_1 = 8'b01111011;
    layers_1_spline_scaler_2 = 8'b11101000;
    layers_1_spline_scaler_3 = 8'b11000000;
    layers_1_spline_scaler_4 = 8'b11111110;
    layers_1_spline_scaler_5 = 8'b10001100;
    layers_1_spline_scaler_6 = 8'b10110011;
    layers_1_spline_scaler_7 = 8'b01000011;
    layers_1_spline_scaler_8 = 8'b00000000;
    layers_1_spline_weight_0 = 8'b01111001;
    layers_1_spline_weight_1 = 8'b01110101;
    layers_1_spline_weight_2 = 8'b01101101;
    layers_1_spline_weight_3 = 8'b10000011;
    layers_1_spline_weight_4 = 8'b01110011;
    layers_1_spline_weight_5 = 8'b01100100;
    layers_1_spline_weight_6 = 8'b10100010;
    layers_1_spline_weight_7 = 8'b10000010;
    layers_1_spline_weight_8 = 8'b01111001;
    layers_1_spline_weight_9 = 8'b01111010;
    layers_1_spline_weight_10 = 8'b01111010;
    layers_1_spline_weight_11 = 8'b01110101;
    layers_1_spline_weight_12 = 8'b01111011;
    layers_1_spline_weight_13 = 8'b01111011;
    layers_1_spline_weight_14 = 8'b01110010;
    layers_1_spline_weight_15 = 8'b01111001;
    layers_1_spline_weight_16 = 8'b01111000;
    layers_1_spline_weight_17 = 8'b01101101;
    layers_1_spline_weight_18 = 8'b01000011;
    layers_1_spline_weight_19 = 8'b01010011;
    layers_1_spline_weight_20 = 8'b10001101;
    layers_1_spline_weight_21 = 8'b01110010;
    layers_1_spline_weight_22 = 8'b11111110;
    layers_1_spline_weight_23 = 8'b10011111;
    layers_1_spline_weight_24 = 8'b01111001;
    layers_1_spline_weight_25 = 8'b01110110;
    layers_1_spline_weight_26 = 8'b01110011;
    layers_1_spline_weight_27 = 8'b10001100;
    layers_1_spline_weight_28 = 8'b10011000;
    layers_1_spline_weight_29 = 8'b10010100;
    layers_1_spline_weight_30 = 8'b10100101;
    layers_1_spline_weight_31 = 8'b10000000;
    layers_1_spline_weight_32 = 8'b01111001;
    layers_1_spline_weight_33 = 8'b01110101;
    layers_1_spline_weight_34 = 8'b01111101;
    layers_1_spline_weight_35 = 8'b10101110;
    layers_1_spline_weight_36 = 8'b10101101;
    layers_1_spline_weight_37 = 8'b10111001;
    layers_1_spline_weight_38 = 8'b10111101;
    layers_1_spline_weight_39 = 8'b01111101;
    layers_1_spline_weight_40 = 8'b01111001;
    layers_1_spline_weight_41 = 8'b01111001;
    layers_1_spline_weight_42 = 8'b01111000;
    layers_1_spline_weight_43 = 8'b01111010;
    layers_1_spline_weight_44 = 8'b10000000;
    layers_1_spline_weight_45 = 8'b01111111;
    layers_1_spline_weight_46 = 8'b01111111;
    layers_1_spline_weight_47 = 8'b01111010;
    layers_1_spline_weight_48 = 8'b01111001;
    layers_1_spline_weight_49 = 8'b01110011;
    layers_1_spline_weight_50 = 8'b01100111;
    layers_1_spline_weight_51 = 8'b10001000;
    layers_1_spline_weight_52 = 8'b01110000;
    layers_1_spline_weight_53 = 8'b01011001;
    layers_1_spline_weight_54 = 8'b10110111;
    layers_1_spline_weight_55 = 8'b10000110;
    layers_1_spline_weight_56 = 8'b01111001;
    layers_1_spline_weight_57 = 8'b01111111;
    layers_1_spline_weight_58 = 8'b10000001;
    layers_1_spline_weight_59 = 8'b01100000;
    layers_1_spline_weight_60 = 8'b10000111;
    layers_1_spline_weight_61 = 8'b10000100;
    layers_1_spline_weight_62 = 8'b01001100;
    layers_1_spline_weight_63 = 8'b01110111;
    layers_1_spline_weight_64 = 8'b01111010;
    layers_1_spline_weight_65 = 8'b10000100;
    layers_1_spline_weight_66 = 8'b10101011;
    layers_1_spline_weight_67 = 8'b10011101;
    layers_1_spline_weight_68 = 8'b01101000;
    layers_1_spline_weight_69 = 8'b10000001;
    layers_1_spline_weight_70 = 8'b00000000;
    layers_1_spline_weight_71 = 8'b01010110;
    layers_2_base_weight_0 = 8'b11111111;
    layers_2_base_weight_1 = 8'b00000000;
    layers_2_base_weight_2 = 8'b10011100;
    layers_2_spline_scaler_0 = 8'b11000111;
    layers_2_spline_scaler_1 = 8'b00000000;
    layers_2_spline_scaler_2 = 8'b11111111;
    layers_2_spline_weight_0 = 8'b10010011;
    layers_2_spline_weight_1 = 8'b10010110;
    layers_2_spline_weight_2 = 8'b10011001;
    layers_2_spline_weight_3 = 8'b10001011;
    layers_2_spline_weight_4 = 8'b10011110;
    layers_2_spline_weight_5 = 8'b10011010;
    layers_2_spline_weight_6 = 8'b01111011;
    layers_2_spline_weight_7 = 8'b10001111;
    layers_2_spline_weight_8 = 8'b01110110;
    layers_2_spline_weight_9 = 8'b00000000;
    layers_2_spline_weight_10 = 8'b11111111;
    layers_2_spline_weight_11 = 8'b11000101;
    layers_2_spline_weight_12 = 8'b01001101;
    layers_2_spline_weight_13 = 8'b10100101;
    layers_2_spline_weight_14 = 8'b10100011;
    layers_2_spline_weight_15 = 8'b10010100;
    layers_2_spline_weight_16 = 8'b10010100;
    layers_2_spline_weight_17 = 8'b10011001;
    layers_2_spline_weight_18 = 8'b10010000;
    layers_2_spline_weight_19 = 8'b10010010;
    layers_2_spline_weight_20 = 8'b10010100;
    layers_2_spline_weight_21 = 8'b10010010;
    layers_2_spline_weight_22 = 8'b10010010;
    layers_2_spline_weight_23 = 8'b10010011;
end


// Layer 0: Input to hidden
assign layer0_out_0 = x1 * layers_0_base_weight_0 + x2 * layers_0_base_weight_1;
assign layer0_out_1 = x1 * layers_0_base_weight_2 + x2 * layers_0_base_weight_3;
assign layer0_out_2 = x1 * layers_0_base_weight_4 + x2 * layers_0_base_weight_5;

// Layer 1: Hidden to hidden
assign layer1_out_0 = layer0_out_0 * layers_1_base_weight_0 + layer0_out_1 * layers_1_base_weight_1 + layer0_out_2 * layers_1_base_weight_2;
assign layer1_out_1 = layer0_out_0 * layers_1_base_weight_3 + layer0_out_1 * layers_1_base_weight_4 + layer0_out_2 * layers_1_base_weight_5;
assign layer1_out_2 = layer0_out_0 * layers_1_base_weight_6 + layer0_out_1 * layers_1_base_weight_7 + layer0_out_2 * layers_1_base_weight_8;

// Layer 2: Hidden to output
assign layer2_out = layer1_out_0 * layers_2_base_weight_0 + layer1_out_1 * layers_2_base_weight_1 + layer1_out_2 * layers_2_base_weight_2;

assign y = layer2_out;

endmodule
